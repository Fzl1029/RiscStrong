///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: Core_Top.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::IGLOO2> <Die::M2GL025> <Package::256 VF>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

//`timescale <time_units> / <precision>

module Core_Top( port1, port2, port3, port4 );
input port1, port2;
output port3;
inout port4;

//<statements>

endmodule

